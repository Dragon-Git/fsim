library rtlLib top.sv,
adder_test.sv,
rtl_adder.sv,
dual_adder.sv;
library gateLib gate_adder.sv;
