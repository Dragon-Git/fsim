library rtlLib rtl_adder.sv,
dual_adder.sv;

library gateLib gate_adder.sv,
gate_adder_alt.sv;

library testLib top.sv,
adder_test.sv;
