library rtlLib rtl_adder.sv;

library gateLib gate_adder.sv,
gate_adder_alt.sv,
dual_adder.sv;

library testLib top.sv,
adder_test.sv;